* jfet model J201 made by https://github.com/dvhx/jfet-model-maker
.model QJ201 NJF(level=2 beta=0.0008163788173493737 delta=0.01 ibd=1.9867767181421779e-13 is=1.4434919873672577e-7 lambda=0.021783763987417805 lfgam=0.0024991991328634977 lfg1=0.000001645567538645927 lfg2=0.0004371620886495023 mvst=0.003385401726772191 mxi=1948.6378263929494 n=30 p=2.303479264306655 q=2.1191771486291744 rd=0.002046721277180671 rs=0.001 vbd=12.43983003685352 vbi=1.1172186177560524 vst=0.15386600309239876 vto=-0.6916396164440355 xi=1752.4527959791917 z=4.968218824272239 acgam=0 cds=0 cgd=0 cgs=0 fc=0.5 hfeta=0 hfe1=0 hfe2=0 hfgam=0 hfg1=0 hfg2=0 taud=0 taug=0 xc=0 af=1 kf=0)
