* jfet model 2N5457
.model Q2N5457 NJF(level=2 beta=0.03313345153507557 delta=5.232699515422614 ibd=1.2561981775200135e-15 is=1.4685541774432905e-10 lambda=0.2781034349079927 lfgam=0.000001 lfg1=0.024299721350373466 lfg2=0.0001179103570268626 mvst=0.7156025730125924 mxi=2.1311996896734335 n=30 p=4.587871842171165 q=2.9221080163665283 rd=0.31201657628420204 rs=0.0010046135746485853 vbd=100 vbi=0.16697844550619542 vst=0.0025416960670707296 vto=-0.24817763851339994 xi=0.09583417695483493 z=100 acgam=0 cds=0 cgd=0 cgs=0 fc=0.5 hfeta=0 hfe1=0 hfe2=0 hfgam=0 hfg1=0 hfg2=0 taud=0 taug=0 xc=0 af=1 kf=0)