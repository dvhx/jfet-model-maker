* jfet model MMBFJ201
.model QMMBFJ201 NJF(level=2 beta=0.000896662032662677 is=3e-12 vto=-0.7942688438190106 delta=0.01 ibd=1.2446786457947927e-15 lambda=0.020523578895410437 lfgam=0.0021458335280504057 lfg1=0.005559062987986806 lfg2=0.0003231192453924478 mvst=0.0000010001509108580035 mxi=153.18973463472332 n=30 p=2.126477686276219 q=2.0772092809108735 rd=0.001 rs=0.0013024536946525222 vbd=56.68319057640032 vbi=9.95066604002855 vst=0.05701116820452227 xi=0.0000010307571946963999 z=1.1391767735628038 acgam=0 cds=0 cgd=0 cgs=0 fc=0.5 hfeta=0 hfe1=0 hfe2=0 hfgam=0 hfg1=0 hfg2=0 taud=0 taug=0 xc=0 af=1 kf=0)