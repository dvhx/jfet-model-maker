* jfet model MMBFJ177LT1G made by https://github.com/dvhx/jfet-model-maker
.model QMMBFJ177LT1G PJF(level=2 beta=0.0019255002930271795 is=3.1754195743859073e-18 vto=-1.2734615523778294 delta=0.39780728413894306 ibd=4.233020763585783e-12 lambda=0.1442323227249739 lfgam=0.0000014773422701272255 lfg1=1e-9 lfg2=0.00009742151122253352 mvst=0.0000018751308248614792 mxi=0.000029975585918661462 n=30 p=7.812707240801008 q=7.42091677526131 rd=64.35027245497552 rs=64.35027245497552 vbd=100 vbi=7.59775994923511 vst=0.0000029890005189806605 xi=0.09925313233382928 z=100 acgam=0 cds=0 cgd=5.5e-9 cgs=1.1e-8 fc=0.5 hfeta=0 hfe1=0 hfe2=0 hfgam=0 hfg1=0 hfg2=0 taud=0 taug=0 xc=0 af=1 kf=0)
