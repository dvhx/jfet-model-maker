* jfet model BF245A
.model QBF245A NJF(level=2 beta=0.03484331174982406 delta=5.402400842072176 ibd=6.096105560585321e-15 is=3.466132230167567e-8 lambda=0.20028254082985852 lfgam=0.000001 lfg1=0.019506023569778545 lfg2=0.000050153069858594216 mvst=0.017529099511278373 mxi=0.000001 n=15.788958660748813 p=4.366468167483658 q=2.8544998771693697 rd=1.5604823102110439 rs=0.0010117014902292344 vbd=71.25331862420573 vbi=0.2510134560172646 vst=0.0000011027201115336583 vto=-0.30274382681557765 xi=7.3949133589070595 z=100 acgam=0 cds=0 cgd=0 cgs=0 fc=0.5 hfeta=0 hfe1=0 hfe2=0 hfgam=0 hfg1=0 hfg2=0 taud=0 taug=0 xc=0 af=1 kf=0)