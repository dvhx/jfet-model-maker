* jfet model TF2123G_E5_AQ3_R
.subckt QTF2123G_E5_AQ3_R_FULL d g s
J_J1 d g s JMOD1
D_D1 s g DMOD1
R_R1 s g 16000000
.model JMOD1 NJF(level=2 beta=0.0015218551373374477 is=3.242812961068422e-12 vto=-0.46211899441556936
  +delta=10.593692303268101 ibd=6.274140933932065e-14 lambda=0.02795532198575133 lfgam=0.0050831513139119
  +lfg1=0.0009883171407377136 lfg2=0.0003885589878250989 mvst=0.5769699295008569 mxi=0.0000015354594023650526
  +n=28.23578450441741 p=2.3485782042625196 q=2.152420967568266 rd=0.20699669276291183 rs=0.03316826991492417
  +vbd=98.70378358277105 vbi=1.429234546265391 vst=0.010494378450143846 xi=1.2478110145177965
  +z=41.471367507655266 acgam=0 cds=0 cgd=0 cgs=0 fc=0.5 hfeta=0 hfe1=0 hfe2=0 hfgam=0 hfg1=0
  +hfg2=0 taud=0 taug=0 xc=0 af=1 kf=0)
.model DMOD1 D(is=1.38738e-10 n=1.73917 rs=0.0043279 cjo=4e-12 vj=0.6 tt=6e-9 m=0.45 bv=100)
.ends
